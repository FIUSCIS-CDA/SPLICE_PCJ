///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SPLICE_PCJ
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: ir25_0 (26-bit), pc31_28 (4-bit)
reg[25:0] ir25_0;
reg[3:0] pc31_28;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: Y (32-bit)
wire[31:0] Y;
///////////////////////////////////////////////////////////////////////////////////

SPLICE_PCJ mySplicer(.ir25_0(ir25_0), .pc31_28(pc31_28), .Y(Y));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: pc31_28=0110, ir25_0=b00001100011000000001101011
$display("Test: pc31_28=0110, ir25_0=b00001100011000000001101011");
pc31_28=4'b0110; ir25_0=26'b00001100011000000001101011;   #10; 
verifyEqual32(Y, {pc31_28, ir25_0, 2'b00});
////////////////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule
